module AND2 (O, I0, I1);
    output O;
    input  I0, I1;

	and A1 (O, I0, I1);

endmodule  
