module AND4 (O, I0, I1, I2, I3);
    output O;
    input  I0, I1, I2, I3;

    and A1 (O, I0, I1, I2, I3);
endmodule