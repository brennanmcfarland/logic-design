module AND3 (O, I0, I1, I2);
    output O;
    input  I0, I1, I2;

    and A1 (O, I0, I1, I2);
endmodule


